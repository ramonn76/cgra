
module branch_selector16x16
(
  input [16-1:0] merge_set_in,
  input [64-1:0] branch_net_conf,
  output [16-1:0] merge_set_out
);

  assign merge_set_out[0] = (branch_net_conf[3:0] == 0 && merge_set_in[0]) | (branch_net_conf[7:4] == 0 && merge_set_in[1]) | (branch_net_conf[11:8] == 0 && merge_set_in[2]) | (branch_net_conf[15:12] == 0 && merge_set_in[3]) | (branch_net_conf[19:16] == 0 && merge_set_in[4]) | (branch_net_conf[23:20] == 0 && merge_set_in[5]) | (branch_net_conf[27:24] == 0 && merge_set_in[6]) | (branch_net_conf[31:28] == 0 && merge_set_in[7]) | (branch_net_conf[35:32] == 0 && merge_set_in[8]) | (branch_net_conf[39:36] == 0 && merge_set_in[9]) | (branch_net_conf[43:40] == 0 && merge_set_in[10]) | (branch_net_conf[47:44] == 0 && merge_set_in[11]) | (branch_net_conf[51:48] == 0 && merge_set_in[12]) | (branch_net_conf[55:52] == 0 && merge_set_in[13]) | (branch_net_conf[59:56] == 0 && merge_set_in[14]) | (branch_net_conf[63:60] == 0 && merge_set_in[15]);
  assign merge_set_out[1] = (branch_net_conf[3:0] == 1 && merge_set_in[0]) | (branch_net_conf[7:4] == 1 && merge_set_in[1]) | (branch_net_conf[11:8] == 1 && merge_set_in[2]) | (branch_net_conf[15:12] == 1 && merge_set_in[3]) | (branch_net_conf[19:16] == 1 && merge_set_in[4]) | (branch_net_conf[23:20] == 1 && merge_set_in[5]) | (branch_net_conf[27:24] == 1 && merge_set_in[6]) | (branch_net_conf[31:28] == 1 && merge_set_in[7]) | (branch_net_conf[35:32] == 1 && merge_set_in[8]) | (branch_net_conf[39:36] == 1 && merge_set_in[9]) | (branch_net_conf[43:40] == 1 && merge_set_in[10]) | (branch_net_conf[47:44] == 1 && merge_set_in[11]) | (branch_net_conf[51:48] == 1 && merge_set_in[12]) | (branch_net_conf[55:52] == 1 && merge_set_in[13]) | (branch_net_conf[59:56] == 1 && merge_set_in[14]) | (branch_net_conf[63:60] == 1 && merge_set_in[15]);
  assign merge_set_out[2] = (branch_net_conf[3:0] == 2 && merge_set_in[0]) | (branch_net_conf[7:4] == 2 && merge_set_in[1]) | (branch_net_conf[11:8] == 2 && merge_set_in[2]) | (branch_net_conf[15:12] == 2 && merge_set_in[3]) | (branch_net_conf[19:16] == 2 && merge_set_in[4]) | (branch_net_conf[23:20] == 2 && merge_set_in[5]) | (branch_net_conf[27:24] == 2 && merge_set_in[6]) | (branch_net_conf[31:28] == 2 && merge_set_in[7]) | (branch_net_conf[35:32] == 2 && merge_set_in[8]) | (branch_net_conf[39:36] == 2 && merge_set_in[9]) | (branch_net_conf[43:40] == 2 && merge_set_in[10]) | (branch_net_conf[47:44] == 2 && merge_set_in[11]) | (branch_net_conf[51:48] == 2 && merge_set_in[12]) | (branch_net_conf[55:52] == 2 && merge_set_in[13]) | (branch_net_conf[59:56] == 2 && merge_set_in[14]) | (branch_net_conf[63:60] == 2 && merge_set_in[15]);
  assign merge_set_out[3] = (branch_net_conf[3:0] == 3 && merge_set_in[0]) | (branch_net_conf[7:4] == 3 && merge_set_in[1]) | (branch_net_conf[11:8] == 3 && merge_set_in[2]) | (branch_net_conf[15:12] == 3 && merge_set_in[3]) | (branch_net_conf[19:16] == 3 && merge_set_in[4]) | (branch_net_conf[23:20] == 3 && merge_set_in[5]) | (branch_net_conf[27:24] == 3 && merge_set_in[6]) | (branch_net_conf[31:28] == 3 && merge_set_in[7]) | (branch_net_conf[35:32] == 3 && merge_set_in[8]) | (branch_net_conf[39:36] == 3 && merge_set_in[9]) | (branch_net_conf[43:40] == 3 && merge_set_in[10]) | (branch_net_conf[47:44] == 3 && merge_set_in[11]) | (branch_net_conf[51:48] == 3 && merge_set_in[12]) | (branch_net_conf[55:52] == 3 && merge_set_in[13]) | (branch_net_conf[59:56] == 3 && merge_set_in[14]) | (branch_net_conf[63:60] == 3 && merge_set_in[15]);
  assign merge_set_out[4] = (branch_net_conf[3:0] == 4 && merge_set_in[0]) | (branch_net_conf[7:4] == 4 && merge_set_in[1]) | (branch_net_conf[11:8] == 4 && merge_set_in[2]) | (branch_net_conf[15:12] == 4 && merge_set_in[3]) | (branch_net_conf[19:16] == 4 && merge_set_in[4]) | (branch_net_conf[23:20] == 4 && merge_set_in[5]) | (branch_net_conf[27:24] == 4 && merge_set_in[6]) | (branch_net_conf[31:28] == 4 && merge_set_in[7]) | (branch_net_conf[35:32] == 4 && merge_set_in[8]) | (branch_net_conf[39:36] == 4 && merge_set_in[9]) | (branch_net_conf[43:40] == 4 && merge_set_in[10]) | (branch_net_conf[47:44] == 4 && merge_set_in[11]) | (branch_net_conf[51:48] == 4 && merge_set_in[12]) | (branch_net_conf[55:52] == 4 && merge_set_in[13]) | (branch_net_conf[59:56] == 4 && merge_set_in[14]) | (branch_net_conf[63:60] == 4 && merge_set_in[15]);
  assign merge_set_out[5] = (branch_net_conf[3:0] == 5 && merge_set_in[0]) | (branch_net_conf[7:4] == 5 && merge_set_in[1]) | (branch_net_conf[11:8] == 5 && merge_set_in[2]) | (branch_net_conf[15:12] == 5 && merge_set_in[3]) | (branch_net_conf[19:16] == 5 && merge_set_in[4]) | (branch_net_conf[23:20] == 5 && merge_set_in[5]) | (branch_net_conf[27:24] == 5 && merge_set_in[6]) | (branch_net_conf[31:28] == 5 && merge_set_in[7]) | (branch_net_conf[35:32] == 5 && merge_set_in[8]) | (branch_net_conf[39:36] == 5 && merge_set_in[9]) | (branch_net_conf[43:40] == 5 && merge_set_in[10]) | (branch_net_conf[47:44] == 5 && merge_set_in[11]) | (branch_net_conf[51:48] == 5 && merge_set_in[12]) | (branch_net_conf[55:52] == 5 && merge_set_in[13]) | (branch_net_conf[59:56] == 5 && merge_set_in[14]) | (branch_net_conf[63:60] == 5 && merge_set_in[15]);
  assign merge_set_out[6] = (branch_net_conf[3:0] == 6 && merge_set_in[0]) | (branch_net_conf[7:4] == 6 && merge_set_in[1]) | (branch_net_conf[11:8] == 6 && merge_set_in[2]) | (branch_net_conf[15:12] == 6 && merge_set_in[3]) | (branch_net_conf[19:16] == 6 && merge_set_in[4]) | (branch_net_conf[23:20] == 6 && merge_set_in[5]) | (branch_net_conf[27:24] == 6 && merge_set_in[6]) | (branch_net_conf[31:28] == 6 && merge_set_in[7]) | (branch_net_conf[35:32] == 6 && merge_set_in[8]) | (branch_net_conf[39:36] == 6 && merge_set_in[9]) | (branch_net_conf[43:40] == 6 && merge_set_in[10]) | (branch_net_conf[47:44] == 6 && merge_set_in[11]) | (branch_net_conf[51:48] == 6 && merge_set_in[12]) | (branch_net_conf[55:52] == 6 && merge_set_in[13]) | (branch_net_conf[59:56] == 6 && merge_set_in[14]) | (branch_net_conf[63:60] == 6 && merge_set_in[15]);
  assign merge_set_out[7] = (branch_net_conf[3:0] == 7 && merge_set_in[0]) | (branch_net_conf[7:4] == 7 && merge_set_in[1]) | (branch_net_conf[11:8] == 7 && merge_set_in[2]) | (branch_net_conf[15:12] == 7 && merge_set_in[3]) | (branch_net_conf[19:16] == 7 && merge_set_in[4]) | (branch_net_conf[23:20] == 7 && merge_set_in[5]) | (branch_net_conf[27:24] == 7 && merge_set_in[6]) | (branch_net_conf[31:28] == 7 && merge_set_in[7]) | (branch_net_conf[35:32] == 7 && merge_set_in[8]) | (branch_net_conf[39:36] == 7 && merge_set_in[9]) | (branch_net_conf[43:40] == 7 && merge_set_in[10]) | (branch_net_conf[47:44] == 7 && merge_set_in[11]) | (branch_net_conf[51:48] == 7 && merge_set_in[12]) | (branch_net_conf[55:52] == 7 && merge_set_in[13]) | (branch_net_conf[59:56] == 7 && merge_set_in[14]) | (branch_net_conf[63:60] == 7 && merge_set_in[15]);
  assign merge_set_out[8] = (branch_net_conf[3:0] == 8 && merge_set_in[0]) | (branch_net_conf[7:4] == 8 && merge_set_in[1]) | (branch_net_conf[11:8] == 8 && merge_set_in[2]) | (branch_net_conf[15:12] == 8 && merge_set_in[3]) | (branch_net_conf[19:16] == 8 && merge_set_in[4]) | (branch_net_conf[23:20] == 8 && merge_set_in[5]) | (branch_net_conf[27:24] == 8 && merge_set_in[6]) | (branch_net_conf[31:28] == 8 && merge_set_in[7]) | (branch_net_conf[35:32] == 8 && merge_set_in[8]) | (branch_net_conf[39:36] == 8 && merge_set_in[9]) | (branch_net_conf[43:40] == 8 && merge_set_in[10]) | (branch_net_conf[47:44] == 8 && merge_set_in[11]) | (branch_net_conf[51:48] == 8 && merge_set_in[12]) | (branch_net_conf[55:52] == 8 && merge_set_in[13]) | (branch_net_conf[59:56] == 8 && merge_set_in[14]) | (branch_net_conf[63:60] == 8 && merge_set_in[15]);
  assign merge_set_out[9] = (branch_net_conf[3:0] == 9 && merge_set_in[0]) | (branch_net_conf[7:4] == 9 && merge_set_in[1]) | (branch_net_conf[11:8] == 9 && merge_set_in[2]) | (branch_net_conf[15:12] == 9 && merge_set_in[3]) | (branch_net_conf[19:16] == 9 && merge_set_in[4]) | (branch_net_conf[23:20] == 9 && merge_set_in[5]) | (branch_net_conf[27:24] == 9 && merge_set_in[6]) | (branch_net_conf[31:28] == 9 && merge_set_in[7]) | (branch_net_conf[35:32] == 9 && merge_set_in[8]) | (branch_net_conf[39:36] == 9 && merge_set_in[9]) | (branch_net_conf[43:40] == 9 && merge_set_in[10]) | (branch_net_conf[47:44] == 9 && merge_set_in[11]) | (branch_net_conf[51:48] == 9 && merge_set_in[12]) | (branch_net_conf[55:52] == 9 && merge_set_in[13]) | (branch_net_conf[59:56] == 9 && merge_set_in[14]) | (branch_net_conf[63:60] == 9 && merge_set_in[15]);
  assign merge_set_out[10] = (branch_net_conf[3:0] == 10 && merge_set_in[0]) | (branch_net_conf[7:4] == 10 && merge_set_in[1]) | (branch_net_conf[11:8] == 10 && merge_set_in[2]) | (branch_net_conf[15:12] == 10 && merge_set_in[3]) | (branch_net_conf[19:16] == 10 && merge_set_in[4]) | (branch_net_conf[23:20] == 10 && merge_set_in[5]) | (branch_net_conf[27:24] == 10 && merge_set_in[6]) | (branch_net_conf[31:28] == 10 && merge_set_in[7]) | (branch_net_conf[35:32] == 10 && merge_set_in[8]) | (branch_net_conf[39:36] == 10 && merge_set_in[9]) | (branch_net_conf[43:40] == 10 && merge_set_in[10]) | (branch_net_conf[47:44] == 10 && merge_set_in[11]) | (branch_net_conf[51:48] == 10 && merge_set_in[12]) | (branch_net_conf[55:52] == 10 && merge_set_in[13]) | (branch_net_conf[59:56] == 10 && merge_set_in[14]) | (branch_net_conf[63:60] == 10 && merge_set_in[15]);
  assign merge_set_out[11] = (branch_net_conf[3:0] == 11 && merge_set_in[0]) | (branch_net_conf[7:4] == 11 && merge_set_in[1]) | (branch_net_conf[11:8] == 11 && merge_set_in[2]) | (branch_net_conf[15:12] == 11 && merge_set_in[3]) | (branch_net_conf[19:16] == 11 && merge_set_in[4]) | (branch_net_conf[23:20] == 11 && merge_set_in[5]) | (branch_net_conf[27:24] == 11 && merge_set_in[6]) | (branch_net_conf[31:28] == 11 && merge_set_in[7]) | (branch_net_conf[35:32] == 11 && merge_set_in[8]) | (branch_net_conf[39:36] == 11 && merge_set_in[9]) | (branch_net_conf[43:40] == 11 && merge_set_in[10]) | (branch_net_conf[47:44] == 11 && merge_set_in[11]) | (branch_net_conf[51:48] == 11 && merge_set_in[12]) | (branch_net_conf[55:52] == 11 && merge_set_in[13]) | (branch_net_conf[59:56] == 11 && merge_set_in[14]) | (branch_net_conf[63:60] == 11 && merge_set_in[15]);
  assign merge_set_out[12] = (branch_net_conf[3:0] == 12 && merge_set_in[0]) | (branch_net_conf[7:4] == 12 && merge_set_in[1]) | (branch_net_conf[11:8] == 12 && merge_set_in[2]) | (branch_net_conf[15:12] == 12 && merge_set_in[3]) | (branch_net_conf[19:16] == 12 && merge_set_in[4]) | (branch_net_conf[23:20] == 12 && merge_set_in[5]) | (branch_net_conf[27:24] == 12 && merge_set_in[6]) | (branch_net_conf[31:28] == 12 && merge_set_in[7]) | (branch_net_conf[35:32] == 12 && merge_set_in[8]) | (branch_net_conf[39:36] == 12 && merge_set_in[9]) | (branch_net_conf[43:40] == 12 && merge_set_in[10]) | (branch_net_conf[47:44] == 12 && merge_set_in[11]) | (branch_net_conf[51:48] == 12 && merge_set_in[12]) | (branch_net_conf[55:52] == 12 && merge_set_in[13]) | (branch_net_conf[59:56] == 12 && merge_set_in[14]) | (branch_net_conf[63:60] == 12 && merge_set_in[15]);
  assign merge_set_out[13] = (branch_net_conf[3:0] == 13 && merge_set_in[0]) | (branch_net_conf[7:4] == 13 && merge_set_in[1]) | (branch_net_conf[11:8] == 13 && merge_set_in[2]) | (branch_net_conf[15:12] == 13 && merge_set_in[3]) | (branch_net_conf[19:16] == 13 && merge_set_in[4]) | (branch_net_conf[23:20] == 13 && merge_set_in[5]) | (branch_net_conf[27:24] == 13 && merge_set_in[6]) | (branch_net_conf[31:28] == 13 && merge_set_in[7]) | (branch_net_conf[35:32] == 13 && merge_set_in[8]) | (branch_net_conf[39:36] == 13 && merge_set_in[9]) | (branch_net_conf[43:40] == 13 && merge_set_in[10]) | (branch_net_conf[47:44] == 13 && merge_set_in[11]) | (branch_net_conf[51:48] == 13 && merge_set_in[12]) | (branch_net_conf[55:52] == 13 && merge_set_in[13]) | (branch_net_conf[59:56] == 13 && merge_set_in[14]) | (branch_net_conf[63:60] == 13 && merge_set_in[15]);
  assign merge_set_out[14] = (branch_net_conf[3:0] == 14 && merge_set_in[0]) | (branch_net_conf[7:4] == 14 && merge_set_in[1]) | (branch_net_conf[11:8] == 14 && merge_set_in[2]) | (branch_net_conf[15:12] == 14 && merge_set_in[3]) | (branch_net_conf[19:16] == 14 && merge_set_in[4]) | (branch_net_conf[23:20] == 14 && merge_set_in[5]) | (branch_net_conf[27:24] == 14 && merge_set_in[6]) | (branch_net_conf[31:28] == 14 && merge_set_in[7]) | (branch_net_conf[35:32] == 14 && merge_set_in[8]) | (branch_net_conf[39:36] == 14 && merge_set_in[9]) | (branch_net_conf[43:40] == 14 && merge_set_in[10]) | (branch_net_conf[47:44] == 14 && merge_set_in[11]) | (branch_net_conf[51:48] == 14 && merge_set_in[12]) | (branch_net_conf[55:52] == 14 && merge_set_in[13]) | (branch_net_conf[59:56] == 14 && merge_set_in[14]) | (branch_net_conf[63:60] == 14 && merge_set_in[15]);
  assign merge_set_out[15] = (branch_net_conf[3:0] == 15 && merge_set_in[0]) | (branch_net_conf[7:4] == 15 && merge_set_in[1]) | (branch_net_conf[11:8] == 15 && merge_set_in[2]) | (branch_net_conf[15:12] == 15 && merge_set_in[3]) | (branch_net_conf[19:16] == 15 && merge_set_in[4]) | (branch_net_conf[23:20] == 15 && merge_set_in[5]) | (branch_net_conf[27:24] == 15 && merge_set_in[6]) | (branch_net_conf[31:28] == 15 && merge_set_in[7]) | (branch_net_conf[35:32] == 15 && merge_set_in[8]) | (branch_net_conf[39:36] == 15 && merge_set_in[9]) | (branch_net_conf[43:40] == 15 && merge_set_in[10]) | (branch_net_conf[47:44] == 15 && merge_set_in[11]) | (branch_net_conf[51:48] == 15 && merge_set_in[12]) | (branch_net_conf[55:52] == 15 && merge_set_in[13]) | (branch_net_conf[59:56] == 15 && merge_set_in[14]) | (branch_net_conf[63:60] == 15 && merge_set_in[15]);

endmodule
